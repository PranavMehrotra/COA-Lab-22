`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date:    16:48:37 10/21/2022 
// Design Name: 
// Module Name:    register_file 
// Project Name: 
// Target Devices: 
// Tool versions: 
// Description: 
//
// Dependencies: 
//
// Revision: 
// Revision 0.01 - File Created
// Additional Comments: 
//
//////////////////////////////////////////////////////////////////////////////////
module register_file(
	input [4:0] rs,
	input [4:0] rt,
	input [4:0] writeReg,
	input [31:0] writeData,
	input clk,
    input rst,
    output reg [31:0] rs_out,
    output reg [31:0] rt_out
    );
    



endmodule
